module main
import lua

fn main() {
	println('Hello Lua!')
}
